library IEEE;
use IEEE.std_logic_1164.all;

-- Declaracion de entidad
entity sum2b_tb is
end;

-- Cuerpo de arquitectura
architecture sum2b_tb_arq of sum2b_tb is
    -- Parte declarativa

	signal a_tb : std_logic_vector(1 downto 0) := "01";
	signal b_tb : std_logic_vector(1 downto 0) := "01";
	signal ci_tb: std_logic := '0';
	signal co_tb: std_logic;
	signal s_tb : std_logic_vector(1 downto 0);
	
begin
    -- Parte descriptiva
	a_tb  <= "11" after 200 ns, "10" after 400 ns;
	b_tb  <= "01" after 300 ns;
	ci_tb <= '1' after 450 ns;
	
	
	sum1b_inst: entity work.sum2b
		port map(
			a_i  => a_tb,
			b_i  => b_tb,
			ci_i => ci_tb,
			s_o  => s_tb,
			co_o => co_tb
			
		);

end;


--
